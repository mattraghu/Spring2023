-- Basic Hello World Program --
